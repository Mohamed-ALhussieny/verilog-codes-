module connection_only(in,out);

parameter width=18;

input  [width-1:0] in;
output [width-1:0] out;

 assign out=in  ;
 endmodule 
